`timescale 1ns/1ns
`include "ebox.svh"

// M8533 CHC
module chc(iCHC CHC);

  // NOTE CHC2,CHC3,CHC4 include Wire-OR of signals by NAME and not
  // directly wired together with lines on the schematic. Beware!

endmodule
