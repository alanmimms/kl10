`timescale 1ns/1ns
// M8521 CHD
module chd(input eboxClk
          );
endmodule // chd
