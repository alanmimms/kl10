`timescale 1ns / 1ps
// M8536 CCL
module ccl(input eboxClk
          /*AUTOARG*/);
endmodule // ccl
