`timescale 1ns/1ns
module cha(input eboxClk
          );
endmodule // cha
