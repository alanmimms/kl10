`timescale 1ns / 1ps
// M8536 CCL
module CCL(input clk
          );
endmodule // CCL
