`ifndef _PI_INTERFACE_
`define _PI_INTERFACE_ 1

interface iPI;
  logic EBUS_CP_GRANT;
  logic EXT_TRAN_REC;
  logic READY;
endinterface

`endif
