`timescale 1ns / 1ps
module PMA(input clk
          );
endmodule // PMA
