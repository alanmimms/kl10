`timescale 1ns / 1ps
// M8533 CHC
module CHC(input clk
          );
endmodule // CHC
