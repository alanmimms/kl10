`timescale 1ns/1ns
`include "ebox.svh"

// M8533 CHC
module chc(iCHC CHC);
endmodule
