// M8520 PAG
module pag(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // pag
