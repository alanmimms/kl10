`timescale 1ns/1ns
// M8531 MBC
module mbc(input eboxClk
          );
endmodule // mbc
