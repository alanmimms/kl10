`timescale 1ns / 1ps
module cha(input eboxClk
          );
endmodule // cha
