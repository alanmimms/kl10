`timescale 1ns / 1ps
// M8521 CHD
module CHD(input clk
          );
endmodule // CHD
