`ifndef _IR_INTERFACE_
`define _IR_INTERFACE_ 1

interface iIR;
  logic ADeq0;
  logic IO_LEGAL;
  logic ADeq0;
  logic ACeq0;
  logic JRST0;
  logic TEST_SATISFIED;
endinterface

`endif
