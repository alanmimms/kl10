`timescale 1ns / 1ps
// M8526 CLK
module CLK(input clk
          );
endmodule // CLK
