`timescale 1ns/1ns
`include "mbox.svh"
module chx(iCHS CHS,
           iMBOX MBOX);

endmodule // chx
