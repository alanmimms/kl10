`timescale 1ns/1ns
// M8536 CCL
module ccl();
endmodule // ccl
