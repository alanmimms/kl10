`ifndef _MBOX_SVH_
 `define _MBOX_SVH_

interface iMBZ;
  logic RD_PSE_WR;
endinterface

`endif
  
    
