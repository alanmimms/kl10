// M8521 CHD
module chd(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // chd
