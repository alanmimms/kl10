`timescale 1ns / 1ps
module CSH(input clk
          );
endmodule // CSH
