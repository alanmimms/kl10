`ifndef _VMA_INTERFACE_
 `define _VMA_INTERFACE_ 1

interface VMA;
  logic [0:35] VMA_HELD_OR_PC;
endinterface

`endif
