`timescale 1ns/1ns
module pma(input eboxClk
          );
endmodule // pma
