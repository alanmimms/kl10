`timescale 1ns / 1ps
// M8520 PAG
module pag(input eboxClk
          );
endmodule // pag
