`timescale 1ns / 1ps
// M8531 MBC
module mbc(input clk
          );
endmodule // mbc
