`timescale 1ns/1ns
module csh();
endmodule // csh
