`timescale 1ns / 1ps
// M8552 DPS
module dps(input clk
          );
endmodule // dps
