`timescale 1ns/1ns
`include "cram-defs.svh"

// M8540 SHM
module shm(input eboxClk,
           iSHM SHM,
           tCRAM CRAM,
           iCON CON,
           iEDP EDP,

           output indexed,
           output ARextended,
           output ARparityOdd
);

endmodule // shm
