`timescale 1ns/1ns
`include "ebox.svh"

// M8542 VMA
module vma(iVMA VMA);

  // XXX temporary
  assign VMA.AC_REF = '0;
endmodule // vma
