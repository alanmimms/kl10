`timescale 1ns / 1ps
// M8537 MBZ
module MBZ(input clk
          );
endmodule // MBZ
