`timescale 1ns/1ns
// M8537 MBZ
module mbz();
endmodule // mbz
