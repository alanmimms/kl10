`timescale 1ns / 1ps
module cha(input clk
          );
endmodule // cha
