`timescale 1ns / 1ps
// M8538 MTR
module mtr(input clk
          );
endmodule // mtr
