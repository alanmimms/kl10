`timescale 1ns / 1ps
// M8542 VMA
module vma(input eboxClk,
           output reg [0:35] VMA_VMAheldOrPC,
           output localACAddress
          /*AUTOARG*/);
endmodule // vma
