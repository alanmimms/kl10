`timescale 1ns / 1ps
// M8531 MBC
module MBC(input clk
          );
endmodule // MBC
