`timescale 1ns / 1ps
module CHA(input clk
          );
endmodule // CHA
