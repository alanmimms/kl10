`timescale 1ns / 1ps
// M8532 PIC
module pic(input eboxClk
          );
endmodule // pic
