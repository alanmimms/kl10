`ifdef TESTBENCH
module kl10pv_tb;
  top kl10pv0();
endmodule
`endif
