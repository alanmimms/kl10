`timescale 1ns / 1ps
// M8533 CHC
module chc(input eboxClk
          );
endmodule // chc
