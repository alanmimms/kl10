`timescale 1ns/1ns
// M8521 CHD
module chd();
endmodule // chd
