`timescale 1ns/1ns
module chx(input eboxClk
          );
endmodule // chx
