// M8525 CON
module con(input eboxClk,
           output loadIR,
           output loadDRAM,
           output longEnable,
           output CON_fmWrite00_17,
           output CON_fmWrite18_35
          /*AUTOARG*/);
  timeunit 1ns;
  timeprecision 1ps;
endmodule // con
