`timescale 1ns / 1ps
// M8525 CON
module con(input eboxClk,
           output loadIR,
           output loadDRAM,
           output longEnable
          /*AUTOARG*/);
endmodule // con
