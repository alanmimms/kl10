`ifndef _SHM_INTERFACE_
`define _SHM_INTERFACE_ 1

interface iSHM;
  logic [0:35] SHM_SH;
  logic [3:0] SHM_XR;
  logic SHM_AR_PAR_ODD;
endinterface

`endif
