// M8536 CCL
module ccl(input eboxClk,
           input eboxReset,
          /*AUTOARG*/);
  timeunit 1ns;
  timeprecision 1ps;
endmodule // ccl
