`timescale 1ns/1ns
// M8542 VMA
module vma(iVMA VMA);

endmodule // vma
