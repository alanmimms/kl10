`timescale 1ns/1ns
`include "ebox.svh"

// M8524 SCD
module scd(iCRAM CRAM,
           iEDP EDP,
           iCTL CTL
);

  iSCD SCD();
endmodule // scd
