`ifndef _APR_INTERFACE_
`define _APR_INTERFACE_ 1

interface iAPR;
  logic [0:2] APR_FMblk;
  logic [0:3] APR_FMadr;
endinterface

`endif
