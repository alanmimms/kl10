`timescale 1ns/1ns
`include "mbox.svh"

// M8537 MBZ
module mbz(iMBZ MBZ);
endmodule // mbz
