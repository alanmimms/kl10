`timescale 1ns/1ns
// M8532 PIC
module pic(input eboxClk
          );
endmodule // pic
