`ifndef 
 `define _PI_INTERFACE_ 1

interface iPI;
  logic GATE_TTL_TO_ECL;
endinterface
`endif
