`timescale 1ns / 1ps
// M8535 CRC
module crc(input eboxClk
          );
endmodule // crc
