module csh(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // csh
