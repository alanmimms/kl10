// M8534 CCW
module ccw(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // ccw

