`timescale 1ns/1ns
// M8542 VMA
module vma(input logic eboxClk,
           input logic eboxReset,
           output logic localACAddress,

           iVMA VMA
);

endmodule // vma
