`timescale 1ns/1ns
`include "cram-defs.svh"
`include "ebus-defs.svh"
// M8524 SCD
module scd(input eboxClk,
           iSCD SCD,
           iCRAM CRAM,
           iEDP EDP,
           iCTL CTL
);

endmodule // scd
