// M8552 DPS
module dps(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // dps
