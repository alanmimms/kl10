`timescale 1ns/1ns
`include "mbox.svh"
module chx(iCSH CSH,
           iMBOX MB);

endmodule // chx
