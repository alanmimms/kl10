module cha(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // cha
