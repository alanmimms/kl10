`timescale 1ns/1ns
`include "ebox.svh"
// M8538 MTR
module mtr();
  iMTR MTR();
endmodule // mtr
