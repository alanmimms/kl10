`timescale 1ns / 1ps
module csh(input eboxClk
          );
endmodule // csh
