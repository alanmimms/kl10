`timescale 1ns/1ns
// M8535 CRC
module crc(input eboxClk
          );
endmodule // crc
