`timescale 1ns/1ns
module chx();
endmodule // chx
