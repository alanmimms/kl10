// M8535 CRC
module crc(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // crc
