// M8537 MBZ
module mbz(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // mbz
