// M8538 MTR
module mtr(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // mtr
