`timescale 1ns / 1ps
module MBOX(input clk,
            input [13:35] vma,
            input vmaACRef,
            input [37:35] mboxGateVMA,
            output [0:35] cacheData,
            input req,
            input read,
            input PSE,
            inputwrite
            );

endmodule // MBOX
