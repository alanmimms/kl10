`ifndef 
 `define _PI_INTERFACE_ 1

interface iPI;
  logic GATE_TTL_TO_ECL;
  logic EBUS_CP_GRANT;
  logic EXT_TRAN_REC;
  logic READY;
endinterface
`endif
