`timescale 1ns / 1ps
module pma(input eboxClk
          );
endmodule // pma
