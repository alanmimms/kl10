`timescale 1ns / 1ps
module csh(input clk
          );
endmodule // csh
