`timescale 1ns/1ns
// M8536 CCL
module ccl(input eboxClk,
           input eboxReset);
endmodule // ccl
