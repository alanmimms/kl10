`timescale 1ns/1ns
// M8537 MBZ
module mbz(input eboxClk
          );
endmodule // mbz
