`timescale 1ns / 1ps
// M8537 MBZ
module mbz(input clk
          );
endmodule // mbz
