`timescale 1ns / 1ps
// M8552 DPS
module DPS(input clk
          );
endmodule // DPS
