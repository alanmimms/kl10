// M8542 VMA
module vma(input eboxClk,
           output reg [0:35] VMA_VMAheldOrPC,
           output localACAddress
          /*AUTOARG*/);
  timeunit 1ns;
  timeprecision 1ps;
endmodule // vma
