`timescale 1ns/1ns
// M8534 CCW
module ccw();
endmodule // ccw

