`timescale 1ns/1ns
// M8538 MTR
module mtr(input eboxClk);
endmodule // mtr
