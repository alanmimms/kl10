`timescale 1ns/1ns
`include "ebox.svh"

// M8542 VMA
module vma(iVMA VMA);
endmodule // vma
