`ifndef _SHM_INTERFACE_
`define _SHM_INTERFACE_ 1

interface iSHM;
  logic [0:35] SH;
  logic [3:0] XR;
  logic AR_PAR_ODD;
endinterface

`endif
