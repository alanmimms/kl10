`timescale 1ns / 1ps
// M8525 CON
module CON(input clk
          );
endmodule // CON
