`timescale 1ns / 1ps
// M8536 CCL
module ccl(input clk
          /*AUTOARG*/);
endmodule // ccl
