`timescale 1ns / 1ps
module chx(input clk
          );
endmodule // chx
