`timescale 1ns / 1ps
// M8532 PIC
module PIC(input clk
          );
endmodule // PIC
