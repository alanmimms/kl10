`timescale 1ns/1ns
// M8520 PAG
module pag();
endmodule // pag
