`ifndef _APR_INTERFACE_
`define _APR_INTERFACE_ 1

interface iAPR;
  logic [0:2] FMblk;
  logic [0:3] FMadr;
endinterface

`endif
