`ifndef _CTL_INTERFACE_
`define _CTL_INTERFACE_ 1

interface iCTL;
  logic CTL_AR00to08_LOAD;
  logic CTL_AR09to17_LOAD;
  logic CTL_ARR_LOAD;
  logic [0:2] CTL_ARL_SEL;
  logic [0:2] CTL_ARR_SEL;
  logic [0:2] CTL_ARXL_SEL;
  logic [0:2] CTL_ARXR_SEL;
  logic CTL_ARX_LOAD;
  logic [0:8] CTL_REG_CTL;
  logic [0:1] CTL_MQ_SEL;
  logic [0:1] CTL_MQM_SEL;
  logic CTL_MQM_EN;
  logic CTL_adToEBUS_L;
  logic CTL_adToEBUS_R;
  logic CTL_DISP_NICOND;
  logic CTL_DISP_RET;
  logic CTL_SPEC_SCM_ALT;
  logic CTL_SPEC_CLR_FPD;
  logic CTL_SPEC_FLAG_CTL;
  logic CTL_SPEC_SP_MEM_CYCLE;
  logic CTL_SPEC_SAVE_FLAGS;
  logic CTL_SPEC_ADX_CRY_36;
  logic CTL_SPEC_GEN_CRY18;
  logic CTL_SPEC_CALL;
  logic CTL_SPEC_SBR_CALL;
  logic CTL_SPEC_XCRY_AR0;
  logic CTL_AD_LONG;
  logic CTL_ADX_CRY_36;
  logic CTL_INH_CRY_18;
  logic CTL_GEN_CRY_18;
  logic CTL_COND_REG_CTL;
  logic CTL_COND_AR_EXP;
  logic CTL_COND_ARR_LOAD;
  logic CTL_COND_ARLR_LOAD;
  logic CTL_COND_ARLL_LOAD;
  logic CTL_COND_AR_CLR;
  logic CTL_COND_ARX_CLR;
  logic CTL_ARL_IND;
  logic [0:1] CTL_ARL_IND_SEL;
  logic CTL_MQ_CLR;
  logic CTL_AR_CLR;
  logic CTL_AR00to11_CLR;
  logic CTL_AR12to17_CLR;
  logic CTL_ARR_CLR;
  logic CTL_ARX_CLR;
  logic CTL_DIAG_CTL_FUNC_00x;
  logic CTL_DIAG_LD_FUNC_04x;
  logic CTL_DIAG_LOAD_FUNC_06x;
  logic CTL_DIAG_LOAD_FUNC_07x;
  logic CTL_DIAG_LOAD_FUNC_072;
  logic CTL_DIAG_LD_FUNC_073;
  logic CTL_DIAG_LD_FUNC_074;
  logic CTL_DIAG_SYNC_FUNC_075;
  logic CTL_DIAG_LD_FUNC_076;
  logic CTL_DIAG_CLK_EDP;
  logic CTL_DIAG_READ_FUNC_11x;
  logic CTL_DIAG_READ_FUNC_12x;
  logic CTL_DIAG_READ_FUNC_13x;
  logic CTL_DIAG_READ_FUNC_14x;
  logic CTL_PI_CYCLE_SAVE_FLAGS;
  logic CTL_LOAD_PC;
  logic CTL_DIAG_STROBE;
  logic CTL_DIAG_READ;
  logic CTL_DIAG_AR_LOAD;
  logic CTL_DIAG_LD_EBUS_REG;
  logic CTL_EBUS_XFER;
  logic CTL_AD_TO_EBUS_L;
  logic CTL_AD_TO_EBUS_R;
  logic CTL_EBUS_T_TO_E_EN;
  logic CTL_EBUS_E_TO_T_EN;
  logic CTL_EBUS_PARITY_OUT;
  logic CTL_DIAG_FORCE_EXTEND;
  logic [0:6] CTL_DIAG_DIAG;
endinterface

`endif
