module chx(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // chx
