`timescale 1ns/1ns
// M8538 MTR
module mtr();
endmodule // mtr
