`timescale 1ns/1ns
module cha();
endmodule // cha
