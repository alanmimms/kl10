`timescale 1ns/1ns
module csh(iCSH CSH);
endmodule // csh
