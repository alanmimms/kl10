`timescale 1ns / 1ps
module pma(input clk
          );
endmodule // pma
