`timescale 1ns / 1ps
// M8521 CHD
module chd(input eboxClk
          );
endmodule // chd
