`timescale 1ns / 1ps
// M8526 CLK
module clk(input clk,
           output mbXfer
          );
endmodule // clk
