// M8531 MBC
module mbc(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // mbc
