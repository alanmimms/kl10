`timescale 1ns / 1ps
// M8542 VMA
module vma(input clk,
           output localACAddress
          /*AUTOARG*/);
endmodule // vma
