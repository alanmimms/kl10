`timescale 1ns/1ns
`include "ebox.svh"

module csh(iAPR APR,
           iCLK CLK,
           iCCL CCL,
           iCSH CSH,
           iMBC MBC,
           iMBX MBX,
           iPMA PMA
           );

  bit clk;
  bit MB_REQ, CHAN_REQ_EN, CYC_TYPE_HOLD, WRITEBACK_T2;
  bit EBOX_REQ_GRANT, EBOX_REQ_EN, NON_EBOX_REQ_GRANT;
  bit CACHE_IDLE_IN_A, CACHE_IDLE_IN_B, CACHE_IDLE_IN_C, CACHE_IDLE_IN_D, CACHE_IDLE_IN_H;
  bit PHASE_CHANGE_COMING, CHAN_RD_T5, E_CACHE_WR_CYC, CACHE_TO_MB_T4;
  bit EBOX_T0, PGRF_CYC, RESET, DATA_DLY_1;
  bit MBOX_RESP, EBOX_RESTART, A_CHANGE_COMING_IN, SBUS_DIAG_3;
  bit ONE_WORD_RD, EBOX_MAP, MAP_PROBLEM, PAGE_FAIL_T2, EBOX_T2;
  bit MB_TEST_PAR_A_IN, LRU_ANY_WR;
  bit PAGE_REFILL_T4_IN, PAGE_REFILL_T4, PAGE_REFILL_T9comma12;
  bit PAGE_REFILL_T10, PAGE_REFILL_T11, PAGE_REFILL_T12, PAGE_REFILL_T13;
  bit EBOX_REFILL_OK, PAGE_REFILL_COMP, PAGE_REFILL_T7;
  bit T0, T1, T2_IN, T3;
  bit CCA_T3, WR_TEST, RD_PSE_2ND_REQ_EN;
  bit e52q3, e52q13, e52q14, e52q15;
  bit EBOX_REQ, CCA_REQ_EN, MB_REQ_GRANT, CACHE_IDLE, EBOX_PAUSE_WRITE, E_CORE_RD_T3;
  bit E_T2_MEM_REF, CCA_CYC_DONE, MEM_BUSY, CHAN_WR_T5, EBOX_RETRY_NEXT;
  bit E_RD_T2_OK, CHAN_T3, WRITEBACK_T1, EBOX_SYNC_HOLD, E_CORE_RD_COMP;
  bit EBOX_READ, E_REQ_EN_CLR, EBOX_RETRY_NEXT_IN;
  bit E_WR_T2, ANY_VALID_MATCH, CACHE_WR_FROM_MEM, RD_FOUND, CACHE_IDLE_IN;
  bit E_WRITEBACK, CORE_BUSY, EBOX_WR_T3, E_RD_T2_CORE_OK, RD_PAUSE_2ND_HALF;
  bit DATA_DLY_2, EBOX_PAUSE, MB_CYC, LOAD_EBUS_REG, EBOX_T3, KI10_PAGING_MODE;
  bit ANY_WRITTEN_MATCH, _0_WD_VAL, _1_WD_VAL, _2_WD_VAL, _3_WD_VAL;
  bit MB_WR_RQ_CLR_NXT, EBOX_TOOK_1_WD, EBOX_T0_IN, WR_DATA_RDY;
  bit PAGE_FAIL_DLY, CSH_T0, EBOX_T1, EBOX_WR_T4, PAGE_FAIL_T3;
  bit EBOX_WR_T4_IN, PAGE_FAIL_HOLD, PAGE_FAIL_DELAY, PAGE_FAIL_HOLD_FF;
  bit DATA_CLR_T2, DATA_CLR_T4, PAGE_REFILL_T8, CHAN_CYC, WR_FROM_MEM_NXT, CCA_CYC;
  bit CHAN_T4, EBOX_SYNC_SEEN, DATA_DLY1, CACHE_WR_IN, WRITE_OK, CCA_INVAL_T4;

  // CSH1 p.24
  always_comb begin
    clk = CLK.CSH;
    CSH.MB_REQ_GRANT = MB_REQ;
    CSH.CHAN_REQ_GRANT = ~MB_REQ & CCL.CHAN_REQ & CHAN_REQ_EN;
    EBOX_REQ_GRANT = ~MB_REQ & CLK.EBOX_REQ & EBOX_REQ_EN & ~CCL.CHAN_REQ;
    CYC_TYPE_HOLD = ~CSH.READY_TO_GO & ~WRITEBACK_T2;

    CSH.EBOX_ERA_GRANT = APR.EBOX_ERA & ~CCL.CHAN_REQ & EBOX_REQ & ~MB_REQ;
    CSH.EBOX_CCA_GRANT = APR.EBOX_CCA & ~CCL.CHAN_REQ & EBOX_REQ & CLK.EBOX_REQ & ~MB_REQ;
    CSH.CCA_REQ_GRANT = MBX.CCA_REQ & ~CCL.CHAN_REQ & CCA_REQ_EN & ~CLK.EBOX_REQ & ~MB_REQ;
    NON_EBOX_REQ_GRANT = PAGE_REFILL_T4 | MB_REQ_GRANT |
                         CSH.CHAN_REQ_GRANT | CSH.CCA_REQ_GRANT;

    CACHE_IDLE_IN_A = PMA.CSH_WRITEBACK_CYC & MBX.CACHE_TO_MB_DONE |
                      ~CSH.READY_TO_GO & CACHE_IDLE |
                      E_CACHE_WR_CYC & CACHE_TO_MB_T4 |
                      CHAN_RD_T5 & PHASE_CHANGE_COMING;

    CACHE_IDLE_IN_B = EBOX_PAUSE_WRITE & E_T2_MEM_REF & PAG.PAGE_OK |
                      (CCA_CYC_DONE | EBOX_WR_T4) |
                      EBOX_T0 & APR.EBOX_LOAD_REG |
                      CACHE_IDLE_IN_C;

    CACHE_IDLE_IN_D = VMA.AC_REF & EBOX_T0 | EBOX_T1 & CLK.EBOX_CYC_ABORT;

    CACHE_IDLE_IN_H = e52q3 | e52q14 | e52q15;

    PGRF_CYC = PMA.PAGE_REFILL_CYC;

    CSH.READY_TO_GO = e52q13 & PAGE_REFILL_T10 |
                      CLK.EBOX_SYNC & CACHE_IDLE |
                      (~CSH.EBOX_CYC | PAGE_REFILL_T4 | RESET) & CACHE_IDLE |
                      ~MCL.VMA_PAUSE & MBOX_RESP & ONE_WORD_RD;

    RESET = CLK.MR_RESET;
  end

  always_ff @(posedge clk) begin
    e52q3 <= CACHE_IDLE_IN_D;
    e52q13 <= ~MEM_BUSY;
    e52q14 <= CACHE_IDLE_IN_A | CHAN_WR_T5 | CACHE_WR_FROM_MEM |
              RESET | CACHE_IDLE_IN_B | EBOX_RETRY_NEXT;
    e52q15 <= CSH.READY_TO_GO & ~EBOX_REQ_GRANT & ~NON_EBOX_REQ_GRANT |
              E_RD_T2_OK & RD_FOUND |
              A_CHANGE_COMING_IN & MBX.SBUS_DIAG_3 |
              CHAN_T3 & ~ANY_VALID_MATCH & CCL.CHAN_TO_MEM;

    CHAN_REQ_EN <= ~WRITEBACK_T1 & ~PAGE_REFILL_T4_IN & ~MEM_BUSY;
    MB_REQ <= MBX.MB_REQ_IN;
    CCA_REQ_EN <= ~WRITEBACK_T1 & ~PAGE_REFILL_T4_IN & ~CORE_BUSY;
  end

  // Note active low symbol
  USR4 e72(.S0('0),
           .D({CSH.EBOX_REQ_GRANT, CSH.MB_REQ_GRANT, CSH.CHAN_REQ_GRANT, CSH.CCA_REQ_GRANT}),
           .S3('0),
           .SEL({2{CYC_TYPE_HOLD}}),
           .Q({CSH.EBOX_CYC, CSH.MB_CYC, CSH.CHAN_CYC, CSH.CCA_CYC}),
           .CLK(clk));


  // CSH2 p.25
  always_comb begin
    CSH.MBOX_RESP_IN = E_RD_T2_OK & RD_FOUND |
                       A_CHANGE_COMING_IN & SBUS_DIAG_3 |
                       ~RESET & (E_CACHE_WR_CYC & CACHE_TO_MB_T4 |
                                 ~EBOX_SYNC_HOLD & DATA_DLY_1 |
                                 MBC.CORE_DATA_VALminus1 & CSH.E_CORE_RD_RQ |
                                 ~E_CORE_RD_COMP & MBOX_RESP & ~EBOX_RESTART) |
                       CACHE_IDLE_IN & CSH.EBOX_CYC;

    EBOX_RESTART = MBOX_RESP & CLK.EBOX_SYNC;
    SBUS_DIAG_3 = MBX.SBUS_DIAG_3;

    E_CACHE_WR_CYC = MCL.VMA_WRITE & CSH.EBOX_CYC & ~EBOX_READ;
    CSH.EBOX_RETRY_REQ = CSH.EBOX_CYC & WRITEBACK_T1 |
                         EBOX_RETRY_NEXT & ~RESET;

    E_REQ_EN_CLR = WRITEBACK_T1 | (E_WRITEBACK & MCL.VMA_READ & PMA.CSH_WRITEBACK_CYC);
    EBOX_RETRY_NEXT_IN = (~MBX.CACHE_BIT | LRU_ANY_WR) &
                         E_WR_T2 & PAG.PAGE_OK & CORE_BUSY &
                         ~ANY_VALID_MATCH |
                         (CSH.ADR_READY &
                          (CORE_BUSY & APR.EBOX_SBUS_DIAG |
                           EBOX_REFILL_OK & PAG.PAGE_REFILL & ~RESET) &
                          CSH.EBOX_CYC) |
                         ~MBC.WRITE_OK & WR_TEST & CSH.EBOX_CYC |
                         ~RD_FOUND & E_RD_T2_OK & CORE_BUSY;
    WR_TEST = CSH.CLEAR_WR_T0 | EBOX_WR_T3;
  end

  always_ff @(posedge clk) begin
    MBOX_RESP <= CSH.MBOX_RESP_IN;

    ONE_WORD_RD <= E_RD_T2_CORE_OK & ~ANY_VALID_MATCH & ~MBX.CACHE_BIT |
                   ~EBOX_RESTART & ONE_WORD_RD & ~CSH.READY_TO_GO;
    RD_PAUSE_2ND_HALF <= ONE_WORD_RD & EBOX_RESTART & EBOX_PAUSE |
                         ~CSH.READY_TO_GO & RD_PAUSE_2ND_HALF;
    RD_PSE_2ND_REQ_EN <= DATA_DLY_2 & RD_PAUSE_2ND_HALF |
                         RD_PSE_2ND_REQ_EN & ~CLK.EBOX_REQ & ~RESET;
    CSH.E_CORE_RD_RQ <= E_RD_T2_CORE_OK & ~RD_FOUND & ANY_VALID_MATCH |
                        ~LRU_ANY_WR & ~ANY_VALID_MATCH | E_RD_T2_CORE_OK |
                        ANY_VALID_MATCH & ~MBX.CACHE_BIT & E_RD_T2_CORE_OK |
                        ~MBC.CORE_DATA_VALID & ~RESET & CSH.E_CORE_RD_RQ;
    EBOX_RETRY_NEXT <= EBOX_RETRY_NEXT_IN;
    EBOX_REQ_EN <= ~CORE_BUSY & ~E_REQ_EN_CLR & ~PAGE_REFILL_T4_IN |
                   MB_CYC & MCL.VMA_READ |
                   RESET |
                   ~E_REQ_EN_CLR & EBOX_REQ_EN & ~EBOX_RETRY_NEXT;
  end


  // CSH3 p.26
  always_comb begin
    LOAD_EBUS_REG = CTL.DIAG_LD_EBUS_REG | PAGE_FAIL_T2 |
                    APR.EBOX_READ_REG & EBOX_T3 & ~MAP_PROBLEM;
    CACHE_IDLE_IN_C = APR.EBOX_READ_REG & EBOX_T3 & ~MAP_PROBLEM | PAGE_FAIL_T3;
    EBOX_MAP = MCL.EBOX_MAP;
    MAP_PROBLEM = MCL.EBOX_MAP &
                  (PAG.PAGE_REFILL | ~KI10_PAGING_MODE) &
                  ~PAG.PAGE_OK;
    CSH.ADR_READY = EBOX_T2 | CSH.T2;
    CSH.ANY_VAL_HOLD_IN = CSH.ADR_READY & ANY_VALID_MATCH |
                          ~CSH.READY_TO_GO & CSH.ANY_VAL_HOLD;
    ANY_WRITTEN_MATCH = CSH._0_VALID_MATCH & CSH._0_ANY_WR |
                        CSH._1_VALID_MATCH & CSH._1_ANY_WR |
                        CSH._2_VALID_MATCH & CSH._2_ANY_WR |
                        CSH._3_VALID_MATCH & CSH._3_ANY_WR;
    RD_FOUND = _0_WD_VAL & CSH._0_VALID_MATCH |
               _1_WD_VAL & CSH._1_VALID_MATCH |
               _2_WD_VAL & CSH._2_VALID_MATCH |
               _3_WD_VAL & CSH._3_VALID_MATCH;
    ANY_VALID_MATCH = CSH._0_VALID_MATCH | CSH._1_VALID_MATCH |
                      CSH._2_VALID_MATCH | CSH._3_VALID_MATCH;
    MB_TEST_PAR_A_IN = DATA_DLY_2 | PAGE_REFILL_T12 | CACHE_WR_FROM_MEM;
    CSH.MATCH_HOLD_IN[0] = (~ANY_VALID_MATCH | CSH._3_VALID_MATCH | CSH._2_VALID_MATCH) &
                           (CSH._2_VALID_MATCH | CSH.LRU_2 | CSH._3_VALID_MATCH);
    CSH.MATCH_HOLD_IN[1] = (~ANY_VALID_MATCH | CSH._3_VALID_MATCH | CSH._1_VALID_MATCH) &
                           (CSH._1_VALID_MATCH | CSH.LRU_1 | CSH._3_VALID_MATCH);
    MB_WR_RQ_CLR_NXT = PAGE_REFILL_T11 | CSH.WR_FROM_MEM_NXT |
                       EBOX_TOOK_1_WD | MBOX.CHAN_READ;
  end

  always_ff @(posedge clk) begin
    CSH.ANY_VAL_HOLD <= CSH.ANY_VAL_HOLD_IN;
    CSH.GATE_VMA_27_33 <= EBOX_T0_IN | (CSH.EBOX_CYC & ~MBX.REFILL_ADR_EN_NXT);
    CSH.ADR_PMA_EN <= ~CSH.EBOX_CYC & ~EBOX_T0_IN & ~MBX.REFILL_ADR_EN_NXT;
  end

  mux2x4 e26(.EN('1),
             .SEL({CSH.LRU_2, CSH.LRU_1}),
             .D0({CSH._0_ANY_WR, CSH._1_ANY_WR, CSH._2_ANY_WR, CSH._3_ANY_WR}),
             .D1(4'b0000),
             .B0(LRU_ANY_WR),
             .B1());


  // CSH4 p.27
  always_comb begin
    CSH.EBOX_T0_IN = CSH.READY_TO_GO & EBOX_REQ_GRANT | CLK.EBOX_REQ & RD_PSE_2ND_REQ_EN;
    E_T2_MEM_REF = ~APR.EBOX_SBUS_DIAG & EBOX_T2 & ~APR.EBOX_READ_REG;
    E_WR_T2 = ~MCL.VMA_PAUSE & E_T2_MEM_REF & ~EBOX_READ;
    E_RD_T2_OK = PAG.PAGE_OK & MCL.VMA_READ & EBOX_T2;
    E_RD_T2_CORE_OK = E_RD_T2_OK & ~CORE_BUSY;
    EBOX_READ = MCL.VMA_READ;
    EBOX_PAUSE_WRITE = ~EBOX_READ & EBOX_PAUSE;
    EBOX_PAUSE = MCL.VMA_PAUSE;
    EBOX_WR_T4_IN = EBOX_WR_T3 & ~EBOX_RETRY_NEXT_IN;
    CSH.REFILL_RAM_WR = APR.EN_REFILL_RAM_WR & EBOX_T2;
  end

  always_ff @(posedge clk) begin
    EBOX_T0 <= CSH.EBOX_T0_IN;
    EBOX_T1 <= EBOX_T0 & ~VMA.AC_REF & ~CACHE_IDLE_IN;
    EBOX_T2 <= EBOX_T1 & ~CLK.EBOX_CYC_ABORT;
    EBOX_T3 <= EBOX_T2;
    CSH.ONE_WORD_WR_T0 <= ~CORE_BUSY & APR.EBOX_SBUS_DIAG & EBOX_T2 |
                          ~MBX.CACHE_BIT & ~ANY_VALID_MATCH & PAG.PAGE_OK &
                          ~CORE_BUSY & ~MCL.VMA_PAUSE & ~EBOX_READ & E_T2_MEM_REF;
    CSH.WRITEBACK_T1 <= ANY_WRITTEN_MATCH & MBX.CSH_CCA_VAL_CORE & CCA_T3 |
                        E_T2_MEM_REF & ~CORE_BUSY & ~EBOX_PAUSE_WRITE &
                        PAG.PAGE_OK & MBX.CACHE_BIT & LRU_ANY_WR & ~ANY_VALID_MATCH;
    WRITEBACK_T2 <= WRITEBACK_T1;

    PAGE_FAIL_DLY <= PAGE_FAIL_HOLD;
    PAGE_FAIL_T2 <= ~(~PAGE_FAIL_DELAY | ~PAGE_FAIL_HOLD);
    PAGE_FAIL_T3 <= PAGE_FAIL_T2;

    DATA_CLR_T2 <= MBC.CSH_DATA_CLR_T3;
    EBOX_WR_T3 <= DATA_CLR_T4 & E_CACHE_WR_CYC |
                  E_WR_T2 & ANY_VALID_MATCH & PAG.PAGE_OK;
    EBOX_WR_T4 <= EBOX_WR_T4_IN;
    CSH.CLEAR_WR_T0 <= PAG.PAGE_OK & ~ANY_VALID_MATCH & E_WR_T2 & MBX.CACHE_BIT & ~LRU_ANY_WR;
    CSH.DATA_CLR_DONE <= MBC.DATA_CLR_DONE_IN & ~CSH.READY_TO_GO |
                         ANY_VALID_MATCH & E_WR_T2 & PAG.PAGE_OK;
  end


  // CSH5 p.28
  always_ff @(posedge clk) begin
    CSH.PAGE_REFILL_T9 <= MBX.CACHE_TO_MB_DONE & PMA.PAGE_REFILL_CYC;
    CSH.PAGE_REFILL_T13 <= PAGE_REFILL_T9comma12;
    PAGE_REFILL_T4 <= PAGE_REFILL_T4_IN;
    PAGE_REFILL_COMP <= PAGE_REFILL_T10 & ~CORE_BUSY |
                        ~EBOX_RESTART & PAGE_REFILL_COMP & ~RESET;
    CSH.PAGE_REFILL_T8 <= PAGE_REFILL_T7;
    PAGE_REFILL_T10 <= CORE_BUSY & ~MBX.MB_SEL_HOLD_FF | PAGE_REFILL_T13;
    PAGE_REFILL_T11 <= PAGE_REFILL_T10;
    CSH.PAGE_REFILL_T12 <= PAGE_REFILL_T11;
    T0 <= ~(~NON_EBOX_REQ_GRANT | ~CSH.READY_TO_GO);
    T1 <= T0;
    CSH.T2 <= T2_IN;
    T3 <= CSH.T2;
    PAGE_REFILL_COMP <= PAGE_REFILL_T10 & ~CORE_BUSY |
                        ~EBOX_RESTART & PAGE_REFILL_COMP & ~RESET;
    PAGE_REFILL_T8 <= PAGE_REFILL_T7;
    CHAN_WR_T5 <= CSH.CHAN_WR_T5_IN;
    CSH.CHAN_T4 <= ANY_VALID_MATCH & CSH.CHAN_T3;
    CSH.CHAN_RD_T5 <= CSH.CHAN_T3 & ~CCL.CHAN_TO_MEM & ~ANY_VALID_MATCH |
                      (MBX.CACHE_TO_MB_DONE & CHAN_CYC & ~RESET &
                       ~CACHE_IDLE_IN & CSH.CHAN_RD_T5);
  end

  always_comb begin
    PAGE_REFILL_T9comma12 = CSH.PAGE_REFILL_T12 & CSH.PAGE_REFILL_T9;
    PAGE_REFILL_T4_IN = ~CORE_BUSY & CSH.EBOX_T3 & EBOX_REFILL_OK & PAG.PAGE_REFILL;
    EBOX_REFILL_OK = (EBOX_MAP | ~APR.EBOX_READ_REG) & ~PAGE_REFILL_COMP;
    PAGE_REFILL_T7 = PAG.PAGE_REFILL_CYC & T3;
    T2_IN = T1 & ~WR_FROM_MEM_NXT;
    CCA_T3 = T3 & CCA_CYC;
    PAGE_REFILL_T7 = PMA.PAGE_REFILL_CYC & T3;
    CSH.CHAN_WR_T5_IN = CCL.CHAN_TO_MEM & CHAN_T4;
    CSH.CHAN_T3 = CHAN_CYC & T3;
  end


  // CSH6 p.29
  always_ff @(posedge clk) begin
    EBOX_SYNC_HOLD <= ~EBOX_T0 & ~RESET & EBOX_SYNC_SEEN;
    CACHE_WR_FROM_MEM <= WR_FROM_MEM_NXT;
    CSH.CHAN_WR_CACHE <= ANY_VALID_MATCH & CCL.CHAN_TO_MEM & CHAN_T3 |
                         CSH.CHAN_WR_CACHE & ~CSH.READY_TO_GO;
    PAGE_FAIL_HOLD_FF <= ~CON.KI10_PAGING_MODE & EBOX_T2 & PAG.PAGE_FAIL |
                         E_T2_MEM_REF & PAG.PAGE_FAIL & ~APR.EBOX_READ_REG |
                         ~CSH.READY_TO_GO & PAGE_FAIL_HOLD_FF & ~APR.EBOX_READ_REG |
                         EBOX_T3 & PAG.PAGE_REFILL & PAGE_REFILL_COMP;
    CSH.PAGE_REFILL_ERROR <= PAGE_REFILL_COMP & PAG.PAGE_REFILL & EBOX_T3 |
                             ~EBOX_RESTART & CSH.PAGE_REFILL_ERROR & ~RESET;
    DATA_DLY_1 <= E_CORE_RD_COMP;
    DATA_DLY_2 <= DATA_DLY1;
    WR_DATA_RDY <= ~ONE_WORD_RD & E_CORE_RD_COMP |
                   WR_DATA_RDY & ~CACHE_WR_IN & ~RESET;
    CSH.CCA_INVAL_T4 <= MBX.CSH_CCA_INVAL_CSH &
                        CCA_T3 &
                        ANY_VALID_MATCH &
                        (~ANY_WRITTEN_MATCH | ~MBX.CSH_CCA_VAL_CORE);
    CSH.CCA_CYC_DONE <= CSH.CCA_INVAL_T4 |
                        ~ANY_VALID_MATCH & CCA_T3 |
                        ~MBX.CSH_CCA_INVAL_CSH & ~ANY_WRITTEN_MATCH & CCA_T3 |
                        ~MBX.CSH_CCA_VAL_CORE & ~MBX.CSH_CCA_INVAL_CSH & CCA_T3;
    CSH.USE_HOLD <= (EBOX_T1 | CSH.USE_HOLD | T2_IN) &
                    ~CSH.READY_TO_GO;
    EBOX_TOOK_1_WD <= EBOX_SYNC_SEEN & ONE_WORD_RD;
  end

  always_comb begin
    EBOX_SYNC_SEEN = EBOX_SYNC_HOLD | EBOX_RESTART;
    WR_FROM_MEM_NXT = EBOX_SYNC_SEEN & WR_DATA_RDY |
                      T1 & MB_CYC & ~RESET;
    CSH.PAGE_FAIL_HOLD = PAGE_FAIL_HOLD_FF;
    E_CORE_RD_COMP = CSH.E_CORE_RD_RQ & MBC.CORE_DATA_VALID;
    CSH.EBOX_LOAD_REG = APR.EBOX_LOAD_REG & EBOX_T0;
    WRITE_OK = MBC.WRITE_OK;
    CSH.CACHE_WR_IN = MBC.CSH_DATA_CLR_T1 & CSH.ONE_WORD_RD & CSH.E_CORE_RD_RQ |
                      EBOX_WR_T3 & WRITE_OK |
                      ~RESET & WR_FROM_MEM_NXT;
    KI10_PAGING_MODE = CON.KI10_PAGING_MODE;
    CSH.MBOX_PT_DIR_WR = ~(~KI10_PAGING_MODE | ~(PAGE_FAIL_T3 | PAGE_REFILL_T12));
    CSH.USE_WR_EN = PAG.PAGE_OK & ANY_VALID_MATCH & EBOX_T2 |
                    ~ONE_WORD_RD & MBC.CSH_DATA_CLR_T2 |
                    MBX.CCA_ALL_PAGES_CYC & CCA_INVAL_T4;
  end


  // CSH7 p.30
  assign CSH.EBUSdriver.driving = CTL.DIAG_READ_FUNC_17x;
  mux e12(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~PAGE_REFILL_COMP, ~CHAN_RD_T5, ~CSH.CHAN_WR_CACHE, ~ONE_WORD_RD,
              ~CSH.E_CORE_RD_RQ, ~CSH.EBOX_RETRY_REQ,
              ~CSH.CCA_INVAL_T4, ~CSH.PAGE_REFILL_ERROR}),
          .q(CSH.EBUSdriver.data[22]));

  mux  e7(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({CSH.CACHE_WR_IN, ~WR_DATA_RDY, ~CSH.CCA_CYC_DONE, ~MBOX_RESP,
              ~CSH.PAGE_FAIL_HOLD, CSH.USE_WR_EN, ~CSH.PAGE_REFILL_T0, ~DATA_DLY_1}),
          .q(CSH.EBUSdriver.data[23]));

  mux e32(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~CSH.MBOX_PT_DIR_WR, ~PAGE_FAIL_T2, ~CSH.CHAN_T4, ~RD_PSE_2ND_REQ_EN,
              ~PAGE_REFILL_T9comma12, ~MB_TEST_PAR_A_IN, ~EBOX_T0, PAGE_FAIL_DLY}),
          .q(CSH.EBUSdriver.data[24]));

  mux  e2(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~WR_TEST, CSH.EBOX_LOAD_REG, CSH.LRU_2, CSH.LRU_1,
              ~CSH._3_ANY_WR, ~CSH._1_ANY_WR, ~CSH._2_ANY_WR, ~CSH._0_ANY_WR}),
          .q(CSH.EBUSdriver.data[25]));

  mux e78(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({CSH.ANY_VAL_HOLD_IN, ~CSH.FILL_CACHE_RD, CSH.READY_TO_GO, ~T1,
              ~CSH_T0, ~T3, ~CSH.T2, ~PAGE_REFILL_T10}),
          .q(CSH.EBUSdriver.data[26]));

  mux e71(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~CSH.DATA_CLR_DONE, ~CHAN_WR_T5, CSH.USE_HOLD, WRITEBACK_T1,
              CSH.ADR_PMA_EN, CSH.GATE_VMA_27_33, CSH.E_CACHE_WR_CYC, CYC_TYPE_HOLD}),
          .q(CSH.EBUSdriver.data[27]));

  mux e73(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~CSH.REFILL_RAM_WR, ~CSH.MB_WR_RQ_CLR_NXT, ~CSH.CCA_CYC, ~CSH.CCA_WRITEBACK,
              ~CSH.EBOX_CYC, ~CSH.MB_CYC, ~CSH.E_WRITEBACK, ~CSH.RD_PAUSE_2ND_HALF}),
          .q(CSH.EBUSdriver.data[28]));

  mux e57(.en(CTL.DIAG_READ_FUNC_17x),
          .sel(CTL.DIAG[4:6]),
          .d({~CSH.EBOX_T3, ~EBOX_T1, ~EBOX_REQ_EN, ~EBOX_T2,
              ~CACHE_IDLE, ~CSH.ONE_WORD_WR_T0, ~CSH.PAGE_REFILL_T4, ~EBOX_WR_T4}),
          .q(CSH.EBUSdriver.data[29]));

  assign E_CORE_RD_T3 = ~EBOX_READ & CSH.EBOX_T3 |
                        EBOX_T3 & CSH.E_CORE_RD_RQ & ~RESET;

  always_ff @(posedge clk) begin
    CSH.FILL_CACHE_RD <= E_CORE_RD_T3 & CSH.E_CORE_RD_RQ |
                         ~EBOX_RESTART & CSH.FILL_CACHE_RD & ~RESET;
    CSH.CCA_WRITEBACK <= WRITEBACK_T1 & CSH.CCA_CYC |
                         ~CACHE_IDLE & CSH.CCA_WRITEBACK;
    CSH.E_WRITEBACK <= WRITEBACK_T1 & CSH.EBOX_CYC |
                       ~E_CORE_RD_T3 & CSH.E_WRITEBACK & ~RESET;
  end
endmodule // csh
