// M8533 CHC
module chc(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // chc
