`timescale 1ns / 1ps
// M8534 CCW
module CCW(input clk
          );
endmodule // CHC
