`timescale 1ns / 1ps
module chx(input eboxClk
          );
endmodule // chx
