`timescale 1ns/1ns
// M8533 CHC
module chc();
endmodule // chc
