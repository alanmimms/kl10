`timescale 1ns/1ns
// M8542 VMA
module vma(input logic eboxClk,
           input logic eboxReset,
           output logic [0:35] VMA_VMAheldOrPC,
           output logic localACAddress);

endmodule // vma
