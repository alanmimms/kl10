`timescale 1ns / 1ps
// M8535 CRC
module CRC(input clk
          );
endmodule // CRC
