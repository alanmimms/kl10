`timescale 1ns/1ns
`include "ebus-defs.svh"
`include "pic.svh"
// M8532 PIC
module pic(input eboxClk,

           iEBUS EBUS,
           tEBUSdriver EBUSdriver,

           iPI PI);

  assign EBUSdriver.driving = 0;       // XXX temporary
endmodule // pic
