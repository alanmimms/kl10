`ifndef _PIC_INTERFACE_
`define _PIC_INTERFACE_ 1

interface iPIC;
  logic PI_EBUS_CP_GRANT;
  logic PI_EXT_TRAN_REC;
  logic PI_READY;
endinterface

`endif
