`timescale 1ns / 1ps
// M8538 MTR
module MTR(input clk
          );
endmodule // MTR
