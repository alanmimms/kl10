`timescale 1ns/1ns
// M8525 CON
module con(input eboxClk,
           output loadIR,
           output loadDRAM,
           output longEnable,
           output CON_fmWrite00_17,
           output CON_fmWrite18_35
          /*AUTOARG*/);
endmodule // con
