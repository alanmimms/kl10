`timescale 1ns/1ns
`include "cram-defs.svh"
`include "ebus-defs.svh"
// M8524 SCD
module scd(iSCD SCD,
           iCRAM CRAM,
           iEDP EDP,
           iCTL CTL
);

endmodule // scd
