`timescale 1ns/1ns
module csh(input eboxClk
          );
endmodule // csh
