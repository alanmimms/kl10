`timescale 1ns/1ns
module pma();
endmodule // pma
