`timescale 1ns / 1ps
module CHX(input clk
          );
endmodule // CHX
