`timescale 1ns / 1ps
// M8520 PAG
module PAG(input clk
          );
endmodule // PAG
