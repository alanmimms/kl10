`timescale 1ns / 1ps
// M8542 VMA
module VMA(input clk
          );
endmodule // VMA
