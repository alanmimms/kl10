`timescale 1ns/1ns
// M8552 DPS
module dps(input eboxClk
          );
endmodule // dps
