`timescale 1ns / 1ps
// M8525 CON
module con(input clk,
           output loadIR,
           output loadDRAM
          );
endmodule // con
