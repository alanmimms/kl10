`timescale 1ns/1ns
`include "ebox.svh"

// M8524 SCD
module scd(iCRAM CRAM,
           iCTL CTL,
           iEDP EDP,
           iSCD SCD
);

endmodule // scd
