// M8532 PIC
module pic(input eboxClk
          );
  timeunit 1ns;
  timeprecision 1ps;
endmodule // pic
