`ifndef _IR_INTERFACE_
`define _IR_INTERFACE_ 1

interface iIR;
  logic IR_ADeq0;
  logic IR_IO_LEGAL;
  logic IR_ACeq0;
  logic IR_JRST0;
  logic IR_TEST_SATISFIED;
endinterface

`endif
